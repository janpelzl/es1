-- simple full adder circuit
entity fa is
    port(
        x: in bit;
        y: in bit;
        cin: in bit;
        s: out bit;
        cout: out bit
    );
end entity;

architecture verhalten of fa is

begin
    s <= (x xor y) xor cin;
    cout <= (x and y) or (x and cin) or (y and cin);

end architecture;
